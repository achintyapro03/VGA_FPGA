module h_sync_controller #(
    parameter front_porch_h = 88,
    parameter sync_width_h  = 44,
    parameter back_porch_h  = 148,
    parameter pixels_h      = 1920
)(
    input clk,
    input reset,
    output reg h_sync,
    output reg video_enable, 
    output reg next_line
);

    reg [11:0] counter;
    wire [11:0] total_pixels;

    assign total_pixels = pixels_h + front_porch_h + sync_width_h + back_porch_h;
    
    always @(posedge clk) begin
        if (reset) begin
            counter <= 12'd0;
            h_sync <= 1'b1;
            video_enable <= 1'b0;
            next_line <= 1'b0;

        end else begin
            if (counter == total_pixels - 1) begin
                counter <= 12'd0;
                next_line <= 1'b1;
            end else begin
                next_line <= 1'b0;
                counter <= counter + 1'b1;
            end

            if (counter < pixels_h) begin
                video_enable <= 1'b1;  
            end else begin
                video_enable <= 1'b0;  
            end

            if (counter >= (pixels_h + front_porch_h) && counter < (pixels_h + front_porch_h + sync_width_h)) begin
                h_sync <= 1'b0;  
            end else begin
                h_sync <= 1'b1;  
            end
        end
    end
endmodule
